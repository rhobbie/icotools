module sim_spiflash (
	input  SPI_FLASH_CS,
	output SPI_FLASH_MISO,
	input  SPI_FLASH_MOSI,
	input  SPI_FLASH_SCLK
);

endmodule
